    -- 0000
    x"02", x"04", x"D4", x"E4", x"90", x"00", x"BC", x"F0",
